`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////
// Company:  NA
// Engineer: Anand J. Roy & Manish Kumar
//
// Create Date:    23:10:06 05/06/20
// Design Name:    
// Module Name:    vending_machine_mod2
// Project Name:   Vending Machine 
// Target Device:  EDGE Spartan 6 FPGA
// Tool versions:  Ise 7.1
// Description:	 Vending machine prototype that dispenses 3 different products of different prices and returns change money according to the money paid.  
//
// Dependencies:	 Actuators that respond to the logic generated by the code.
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////
module vending_machine_mod2(delivered,change,cancel,item_number,i,j,rst,clk);
input cancel,i,j,rst,clk;
input [1:0]item_number;
output reg delivered,change;
reg [2:0] state, NS;
parameter  s0=3'b000,s1=3'b001,s2=3'b010,s3=3'b011,s4=3'b100,s5=3'b101,s6=3'b110,s7=3'b111;

always @ (posedge clk or negedge rst)
if (~rst) 
	state=s0;
else 
	state = NS;

always @ (state or i or j or cancel or item_number)
case(item_number)

	2'b11: // Product C - Cost Rs.3
	begin
		case(state)
		s0: NS = cancel?s0:(i?(j?s2:s1):s0);
		s1: NS = cancel?s5:(i?(j?s3:s2):s1);
		s2: NS = cancel?s6:(i?(j?s4:s3):s2);
		s3: NS = s0;
		s4: NS = s0;
		s5: NS = s0;
		s6: NS = s5;
		endcase

		assign {delivered,change} = {(state[0] & state[1] & ~state[2])|(~state[0] & ~state[1] & state[2]),(state[2] & ~state[1])|(state[2] & ~state[0])};
	end
	2'b10: // Product B - Cost Rs.2
	begin
		case(state)
		s0: NS = cancel?s0:(i?(j?s2:s1):s0);
		s1: NS = cancel?s4:(i?(j?s3:s2):s1);
		s2: NS = s0;
		s3: NS = s0;
		s4: NS = s0;
		endcase
		
		assign {delivered,change} = {(state[1] & ~state[2]),(~state[0] & ~state[1] & state[2])|(state[0] & state[1] & ~state[2])};
	end
	2'b01: // Product A - Cost Re.1
	begin
		case(state)
		s0: NS = cancel?s0:(i?(j?s2:s1):s0);
		s1: NS = s0;
		s2: NS = s0;
		endcase
		
		assign {delivered,change} = {((state[0] & ~state[1] & ~state[2])|(~state[0] & state[1] & ~state[2])),(~state[0] & state[1] & ~state[2])};
	end
	endcase	
		
endmodule